module ExampleModule #(
    parameter WIDTH = 8,
    parameter DEPTH = 16,
    parameter ADDR_WIDTH = 4
)(
    // Inputs
    input wire clk,
    input wire reset,
    input wire [WIDTH-1:0] data_in,
    input logic [DEPTH-1:0] enable,
    input bit [7:0] config,
    input reg [3:0] mode,
    input wire [15:0] address,
    input [31:0] instruction,
    input wire start,
    input wire [ADDR_WIDTH-1:0] write_addr,
    input logic [15:0] mask,
    input wire init,
    input bit stop,
    input [WIDTH-1:0] threshold,
    input logic [3:0] status,
    input wire ready,
    input bit [7:0] flag,
    input reg [DEPTH-1:0] counter,
    input logic [WIDTH-1:0] buffer,
    input wire [WIDTH-1:0] temp,
    input bit [3:0] cmd,
    input reg [7:0] control,
    input wire [15:0] shift,
    input logic [7:0] interrupt,
    input wire done,
    input [WIDTH-1:0] data_in_ext,

    // Outputs
    output wire [WIDTH-1:0] data_out,
    output logic [DEPTH-1:0] status_out,
    output bit [7:0] config_out,
    output reg [3:0] mode_out,
    output wire [15:0] address_out,
    output [31:0] result,
    output wire complete,
    output wire [ADDR_WIDTH-1:0] read_addr,
    output logic [15:0] mask_out,
    output wire init_done,
    output bit stop_ack,
    output [WIDTH-1:0] threshold_out,
    output logic [3:0] status_flag,
    output wire ready_signal,
    output bit [7:0] error_flag,
    output reg [DEPTH-1:0] counter_out,
    output logic [WIDTH-1:0] buffer_out,
    output wire [WIDTH-1:0] temp_out,
    output bit [3:0] cmd_out,
    output reg [7:0] control_out,
    output wire [15:0] shift_out,
    output logic [7:0] interrupt_out,
    output wire task_done,
    output [WIDTH-1:0] data_out_ext,

    // Inouts
    inout wire [WIDTH-1:0] bidir_data,
    inout logic [DEPTH-1:0] bidir_status,
    inout bit [7:0] bidir_config,
    inout reg [3:0] bidir_mode,
    inout wire [15:0] bidir_address,
    inout [31:0] bidir_instruction,
    inout wire bidir_start,
    inout wire [ADDR_WIDTH-1:0] bidir_write_addr,
    inout logic [15:0] bidir_mask,
    inout wire bidir_init,
    inout bit bidir_stop
);

// Module implementation here

endmodule
