--doc init
--This is module NO8
--inputs:
--a : input 1
--outputs:
--b : output 1
--doc end