--doc init
--This is module NO6
--inputs:
--a : input 1
--outputs:
--b : output 1
--doc end